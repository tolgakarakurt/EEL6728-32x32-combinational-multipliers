------------------------------------------------------------------------------------------
--Karakurt--------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.all;
------------------------------------------------------------------------------------------
entity vmul32x32i is
	port (
		X: in UNSIGNED (31 downto 0);
		Y: in UNSIGNED (31 downto 0);
		P: out UNSIGNED (63 downto 0)
		);
end vmul32x32i;
------------------------------------------------------------------------------------------
architecture vmul32x32i_arch of vmul32x32i is
begin
	P <= X * Y;
end vmul32x32i_arch;
------------------------------------------------------------------------------------------
