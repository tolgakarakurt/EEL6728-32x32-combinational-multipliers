------------------------------------------------------------------------------------------
--Karakurt--------------------------------------------------------------------------------
------------------------------------------------------------------------------------------
 ---------------------------------------
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;
 ---------------------------------------
 ENTITY AND2 IS
	--GENERIC(delay: time :=111 ps);
 	port( I0, I1: in STD_LOGIC;
		   O: out STD_LOGIC );
 END AND2;
 ---------------------------------------
 ARCHITECTURE and2_arch OF AND2 IS
 BEGIN
	O <= I0 AND I1; --AFTER delay;
 END ARCHITECTURE;
 ---------------------------------------
